`timescale 1 ns / 1 ps
module fifomem_TB #(parameter WORDSIZE = 8,
                parameter ADDRSIZE = 8)
              ();
endmodule